module register12_r_en(q, clk, reset_n, en, d);	//12-bits reset_n / en register
	input clk, reset_n, en;
	input [11:0] d;
	output reg [11:0] q;
	
	always@(posedge clk or negedge reset_n)		//Operate when clk and reset_n is changed
	begin
		if(reset_n == 0)		q <= 12'b0;			//reset
		else if(en)				q <= d;				//store
		else						q <= q;				//write
	end
endmodule
